
// Accurate Multiplier


module accumul(
    input [1:0] a,
    input [1:0] b,
    output [3:0] out
);

    assign out = a * b;

endmodule